module ALU( 
	input	[31:0]	a,
	input	[31:0]	b,
	input	[3:0]	aluop,
	output	[31:0]	result,
	output			zero
);

	wire [31:0]	logicout;	// output of the logic block
	wire [31:0]	addout;		// adder subtractor out
	wire [31:0]	arithout;	// output after alt
	wire [31:0]	n_b;		// inverted b
	wire [31:0]	sel_b;		// select b or n_b;
	wire [31:0]	slt;		// output of the slt extension

	wire [1:0]	logicsel;	// lower two bits of aluop;

	// logic select 
	assign logicsel =	aluop[1:0];
	assign logicout =	(logicsel == 2'b00) ? a & b :
						(logicsel == 2'b01) ? a | b :
						(logicsel == 2'b10) ? a ^ b :
											~(a | b);

	// adder subtractor
	assign n_b = ~b;  // invert b
	assign sel_b = (aluop[1]) ? n_b : b ;
	assign addout = a + sel_b + aluop[1];

	// set less than operator
	assign slt = {31'b0, addout[31]};
	
	// arith out
	assign arithout = (aluop[3]) ? slt : addout;
	
	// final out
	assign result = (aluop[2]) ? logicout : arithout;
	// the zero
	assign zero = (result == 32'b0) ? 1 : 0;

endmodule
