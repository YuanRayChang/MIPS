module InstructionMemory(
	input	[5:0]	A,	// Address of the Instruction max 64 instructions
	output	[31:0]	RD	// Value at Address
);

	reg [31:0] InsArr [63:0];	// Array holding the memory 64 entries each 32 bits

	initial
	begin
		// Initialize the array with this content
		$readmemh("insmem_direction_h.txt", InsArr);
	end

	assign RD = InsArr[A];   // The Read Data (RD) output corresponds to the Address (A)

endmodule